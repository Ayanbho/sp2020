
/* 
Copyright (c) 2019, IIT Madras All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.  
* Redistributions in binary form must reproduce the above copyright notice, this list of 
  conditions and the following disclaimer in the documentation and/or other materials provided 
  with the distribution.  
* Neither the name of IIT Madras  nor the names of its contributors may be used to endorse or 
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT 
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------

This file has been generated by ProtoSynth.
Time of Generation: 2020-01-23 18:18:07.528693

*/

package coherence_types;

`include "coherence.defines"

typedef enum { 
  Load,
  Store,
  Evict,
  None
} Access deriving (Eq, Bits, FShow);


typedef enum { 
  GetS,
  GetS_Ack,
  GetM,
  GetM_Ack_D,
  GetM_Ack_AD,
  Inv_Ack,
  Upgrade,
  PutS,
  Put_Ack,
  WB,
  PutM,
  Inv,
  Fwd_GetS,
  Fwd_GetM
} MessageType deriving (Eq, Bits, FShow);


typedef enum { 
  Cacheline_state_I,
  Cacheline_state_I_Load,
  Cacheline_state_I_Store,
  Cacheline_state_I_Store_GetM_Ack_AD,
  Cacheline_state_M,
  Cacheline_state_M_Evict,
  Cacheline_state_M_Evict_Fwd_GetM,
  Cacheline_state_S,
  Cacheline_state_S_Evict,
  Cacheline_state_S_Store,
  Cacheline_state_S_Store_GetM_Ack_AD
} Cacheline_state deriving (Eq, Bits, FShow);


typedef enum { 
  Dict_I,
  Dict_M,
  Dict_M_GetS,
  Dict_S
} Dict deriving (Eq, Bits, FShow);



typedef union tagged {
 
  Bit#(TLog#(`NrCaches)) Caches;
  void Directory;
} Machines deriving(Eq, Bits, FShow);

typedef struct {
  Bit#(a) address;
  MessageType msgtype;
  Machines src;
  Machines dst;
  Bit#(TLog#(`NrCaches)) acksExpected;
  Bit#(TMul#(8,w)) cl;

} Message #(numeric type a, numeric type w) deriving(Eq, Bits, FShow);

typedef struct {
  Cacheline_state state;
  Access perm;
  Bit#(TMul#(8,w)) cl;
  Bit#(TLog#(`NrCaches)) acksReceived;
  Bit#(TLog#(`NrCaches)) acksExpected;
  Machines id;

} ENTRY_Cacheline_state #(numeric type w) deriving(Eq, Bits, FShow);


typedef struct {
    Bool stall;
    ENTRY_Cacheline_state#(w) new_cle;
    Maybe#( Message#(a,w) ) send_resp1;
    Maybe#( Message#(a,w) ) send_resp2;
} Cacheline_stateReturn #(numeric type a, numeric type w) deriving(Bits, Eq, FShow);


typedef struct {
  Dict state;
  Access perm;
  Bit#(TMul#(8,w)) cl;
  V_NrCaches_OBJSET_sv sv;
  Machines owner;
  Machines id;

} ENTRY_Dict #(numeric type w) deriving(Eq, Bits, FShow);


typedef struct {
    Bool stall;
    ENTRY_Dict#(w) new_cle;
    Maybe#( Message#(a,w) ) send_resp1;
    Maybe#( Message#(a,w) ) send_fwd1;
    Maybe#(Tuple2#(Message#(a,w),Bit#(`NrCaches))) send_multicast;
} DictReturn #(numeric type a, numeric type w) deriving(Bits, Eq, FShow);

typedef Bit#(`NrCaches) V_NrCaches_OBJSET_sv;
typedef Bit#(TLog#(`NrCaches)) Cnt_V_NrCaches_OBJSET_sv;


function Message#(a,w) fn_Request(Bit#(a) address, MessageType msgtype, Machines src, Machines dst);
  Message#(a,w) msg;
  msg.address = address;
  msg.msgtype = msgtype;
  msg.src = src;
  msg.dst = dst;
  msg.acksExpected = ?;
  msg.cl = ?;
  return msg;
endfunction

function Message#(a,w) fn_Ack(Bit#(a) address, MessageType msgtype, Machines src, Machines dst);
  Message#(a,w) msg;
  msg.address = address;
  msg.msgtype = msgtype;
  msg.src = src;
  msg.dst = dst;
  msg.acksExpected = ?;
  msg.cl = ?;
  return msg;
endfunction

function Message#(a,w) fn_Resp(Bit#(a) address, MessageType msgtype, Machines src, Machines dst, Bit#(TMul#(8,w)) cl);
  Message#(a,w) msg;
  msg.address = address;
  msg.msgtype = msgtype;
  msg.src = src;
  msg.dst = dst;
  msg.acksExpected = ?;
  msg.cl = cl;
  return msg;
endfunction

function Message#(a,w) fn_RespAck(Bit#(a) address, MessageType msgtype, Machines src, Machines dst, Bit#(TMul#(8,w)) cl, Bit#(TLog#(`NrCaches)) acksExpected);
  Message#(a,w) msg;
  msg.address = address;
  msg.msgtype = msgtype;
  msg.src = src;
  msg.dst = dst;
  msg.acksExpected = acksExpected;
  msg.cl = cl;
  return msg;
endfunction



function V_NrCaches_OBJSET_sv fn_Clear(V_NrCaches_OBJSET_sv sv);
  return 0;
endfunction

function V_NrCaches_OBJSET_sv fn_RemoveElement(V_NrCaches_OBJSET_sv sv, Machines src);
  if ( src matches tagged Caches .c)
    sv[c] = 0;
  return sv;
endfunction

function V_NrCaches_OBJSET_sv fn_AddElement(V_NrCaches_OBJSET_sv sv, Machines src);
  if ( src matches tagged Caches .c)
      sv[c] = 1;
  return sv;
endfunction

function Bool fn_IsElement (V_NrCaches_OBJSET_sv sv, Machines i);
  if ( i matches tagged Caches .c)
    return unpack(sv[c]);
  else
    return False;
endfunction

function Cnt_V_NrCaches_OBJSET_sv fn_VectorCount (V_NrCaches_OBJSET_sv sv);
  return truncate(pack(countOnes(sv)));
endfunction




function Cacheline_stateReturn#(a,w) func_Cacheline_state(Message#(a,w) inmsg, ENTRY_Cacheline_state#(w) cle);
  Message#(a,w) msg; 
  let address = inmsg.address ;
  Bool stall = False;
  Maybe#(Message#(a,w)) send_resp1 = tagged Invalid;
  Maybe#(Message#(a,w)) send_resp2 = tagged Invalid;
  Maybe#(Message#(a,w)) enq_defermsg1 = tagged Invalid;
  Maybe#(Message#(a,w)) enq_defermsg2 = tagged Invalid;
  Bool send_defermsg = False;
  case (cle.state) 

    Cacheline_state_I: begin
    case (inmsg.msgtype)
       default: stall = True;
    endcase
    end

    Cacheline_state_I_Load: begin
    case (inmsg.msgtype)
      GetS_Ack: begin
        cle.cl = inmsg.cl;
        cle.state = Cacheline_state_S;
        cle.perm = Load;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_I_Store: begin
    case (inmsg.msgtype)
      GetM_Ack_AD: begin
        cle.acksExpected = inmsg.acksExpected;
        cle.cl = inmsg.cl;
        if (cle.acksExpected == cle.acksReceived) begin
        cle.state = Cacheline_state_M;
        cle.perm = Store;

      end

        else begin
        cle.state = Cacheline_state_I_Store_GetM_Ack_AD;
        cle.perm = None;
        end

      end

      GetM_Ack_D: begin
        cle.cl = inmsg.cl;
        cle.state = Cacheline_state_M;
        cle.perm = Store;

      end

      Inv_Ack: begin
        cle.acksReceived = cle.acksReceived+1;
        cle.state = Cacheline_state_I_Store;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_I_Store_GetM_Ack_AD: begin
    case (inmsg.msgtype)
      Inv_Ack: begin
        cle.acksReceived = cle.acksReceived+1;
        if (cle.acksExpected == cle.acksReceived) begin
        cle.state = Cacheline_state_M;
        cle.perm = Store;

      end

        else begin
        cle.state = Cacheline_state_I_Store_GetM_Ack_AD;
        cle.perm = None;
        end

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_M: begin
    case (inmsg.msgtype)
      Fwd_GetM: begin
        msg = fn_Resp(address,GetM_Ack_D,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Cacheline_state_I;
        cle.perm = None;

      end

      Fwd_GetS: begin
        msg = fn_Resp(address,GetS_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        msg = fn_Resp(address,WB,cle.id,tagged Directory,cle.cl);
        send_resp2 = tagged Valid msg;
        cle.state = Cacheline_state_S;
        cle.perm = Load;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_M_Evict: begin
    case (inmsg.msgtype)
      Fwd_GetM: begin
        msg = fn_Resp(address,GetM_Ack_D,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Cacheline_state_M_Evict_Fwd_GetM;
        cle.perm = None;

      end

      Fwd_GetS: begin
        msg = fn_Resp(address,GetS_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        msg = fn_Resp(address,WB,cle.id,tagged Directory,cle.cl);
        send_resp2 = tagged Valid msg;
        cle.state = Cacheline_state_S_Evict;
        cle.perm = None;

      end

      Put_Ack: begin
        cle.state = Cacheline_state_I;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_M_Evict_Fwd_GetM: begin
    case (inmsg.msgtype)
      Put_Ack: begin
        cle.state = Cacheline_state_I;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_S: begin
    case (inmsg.msgtype)
      Inv: begin
        msg = fn_Resp(address,Inv_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Cacheline_state_I;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_S_Evict: begin
    case (inmsg.msgtype)
      Inv: begin
        msg = fn_Resp(address,Inv_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Cacheline_state_M_Evict_Fwd_GetM;
        cle.perm = None;

      end

      Put_Ack: begin
        cle.state = Cacheline_state_I;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_S_Store: begin
    case (inmsg.msgtype)
      GetM_Ack_AD: begin
        cle.acksExpected = inmsg.acksExpected;
        if (cle.acksExpected == cle.acksReceived) begin
        cle.state = Cacheline_state_M;
        cle.perm = Store;

      end

        else begin
        cle.state = Cacheline_state_S_Store_GetM_Ack_AD;
        cle.perm = Load;
        end

      end

      GetM_Ack_D: begin
        cle.state = Cacheline_state_M;
        cle.perm = Store;

      end

      Inv: begin
        msg = fn_Resp(address,Inv_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Cacheline_state_I_Store;
        cle.perm = None;

      end

      Inv_Ack: begin
        cle.acksReceived = cle.acksReceived+1;
        cle.state = Cacheline_state_S_Store;
        cle.perm = Load;

      end

       default: stall = True;
    endcase
    end

    Cacheline_state_S_Store_GetM_Ack_AD: begin
    case (inmsg.msgtype)
      Inv_Ack: begin
        cle.acksReceived = cle.acksReceived+1;
        if (cle.acksExpected == cle.acksReceived) begin
        cle.state = Cacheline_state_M;
        cle.perm = Store;

      end

        else begin
        cle.state = Cacheline_state_S_Store_GetM_Ack_AD;
        cle.perm = Load;
        end

      end

       default: stall = True;
    endcase
    end

endcase
return Cacheline_stateReturn { stall : stall, new_cle: cle, send_resp1: send_resp1, send_resp2: send_resp2};
endfunction
function DictReturn#(a,w) func_Dict(Message#(a,w) inmsg, ENTRY_Dict#(w) cle);
  Message#(a,w) msg; 
  Bool stall = False;
  let address = inmsg.address ;
  Maybe#(Message#(a,w)) send_resp1 = tagged Invalid;
  Maybe#(Message#(a,w)) send_fwd1 = tagged Invalid;
  Maybe#(Tuple2#(Message#(a,w),Bit#(`NrCaches))) send_multicast = tagged Invalid;
  case (cle.state) 

    Dict_I: begin
    case (inmsg.msgtype)
      GetM: begin
        msg = fn_RespAck(address,GetM_Ack_AD,cle.id,inmsg.src,cle.cl,fn_VectorCount (cle.sv));
        send_resp1 = tagged Valid msg;
        cle.owner = inmsg.src;
        cle.state = Dict_M;
        cle.perm = None;

      end

      GetS: begin
        cle.sv = fn_AddElement(cle.sv,inmsg.src);
        msg = fn_Resp(address,GetS_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Dict_S;
        cle.perm = None;

      end

      PutM: begin
        msg = fn_Ack(address,Put_Ack,cle.id,inmsg.src);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        if (cle.owner == inmsg.src) begin
        cle.cl = inmsg.cl;
        cle.state = Dict_I;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_I;
        cle.perm = None;
        end

      end

      PutS: begin
        msg = fn_Resp(address,Put_Ack,cle.id,inmsg.src,cle.cl);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        if (fn_VectorCount (cle.sv) == 0) begin
        cle.state = Dict_I;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_I;
        cle.perm = None;
        end

      end

      Upgrade: begin
        msg = fn_RespAck(address,GetM_Ack_AD,cle.id,inmsg.src,cle.cl,fn_VectorCount (cle.sv));
        send_resp1 = tagged Valid msg;
        cle.owner = inmsg.src;
        cle.state = Dict_M;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Dict_M: begin
    case (inmsg.msgtype)
      GetM: begin
        msg = fn_Request(address,Fwd_GetM,inmsg.src,cle.owner);
        send_fwd1 = tagged Valid msg;
        cle.owner = inmsg.src;
        cle.state = Dict_M;
        cle.perm = None;

      end

      GetS: begin
        msg = fn_Request(address,Fwd_GetS,inmsg.src,cle.owner);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_AddElement(cle.sv,inmsg.src);
        cle.sv = fn_AddElement(cle.sv,cle.owner);
        cle.state = Dict_M_GetS;
        cle.perm = None;

      end

      PutM: begin
        msg = fn_Ack(address,Put_Ack,cle.id,inmsg.src);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        if (cle.owner == inmsg.src) begin
        cle.cl = inmsg.cl;
        cle.state = Dict_I;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_M;
        cle.perm = None;
        end

      end

      PutS: begin
        msg = fn_Resp(address,Put_Ack,cle.id,inmsg.src,cle.cl);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        if (fn_VectorCount (cle.sv) == 0) begin
        cle.state = Dict_M;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_M;
        cle.perm = None;
        end

      end

      Upgrade: begin
        msg = fn_Request(address,Fwd_GetM,inmsg.src,cle.owner);
        send_fwd1 = tagged Valid msg;
        cle.owner = inmsg.src;
        cle.state = Dict_M;
        cle.perm = None;

      end

       default: stall = True;
    endcase
    end

    Dict_M_GetS: begin
    case (inmsg.msgtype)
      WB: begin
        if (inmsg.src == cle.owner) begin
        cle.cl = inmsg.cl;
        cle.state = Dict_S;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_M_GetS;
        cle.perm = None;
        end

      end

       default: stall = True;
    endcase
    end

    Dict_S: begin
    case (inmsg.msgtype)
      GetM: begin
        if (fn_IsElement (cle.sv,inmsg.src)) begin
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        msg = fn_RespAck(address,GetM_Ack_AD,cle.id,inmsg.src,cle.cl,fn_VectorCount (cle.sv));
        send_resp1 = tagged Valid msg;
        cle.state = Dict_M;
        cle.perm = None;
        msg = fn_Ack(address,Inv,inmsg.src,inmsg.src);
        send_multicast = tagged Valid tuple2(msg,cle.sv);
        cle.owner = inmsg.src;
        cle.sv = fn_Clear(cle.sv);

      end

        else begin
        msg = fn_RespAck(address,GetM_Ack_AD,cle.id,inmsg.src,cle.cl,fn_VectorCount (cle.sv));
        send_resp1 = tagged Valid msg;
        cle.state = Dict_M;
        cle.perm = None;
        msg = fn_Ack(address,Inv,inmsg.src,inmsg.src);
        send_multicast = tagged Valid tuple2(msg,cle.sv);
        cle.owner = inmsg.src;
        cle.sv = fn_Clear(cle.sv);
        end

      end

      GetS: begin
        cle.sv = fn_AddElement(cle.sv,inmsg.src);
        msg = fn_Resp(address,GetS_Ack,cle.id,inmsg.src,cle.cl);
        send_resp1 = tagged Valid msg;
        cle.state = Dict_S;
        cle.perm = None;

      end

      PutM: begin
        msg = fn_Ack(address,Put_Ack,cle.id,inmsg.src);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        if (cle.owner == inmsg.src) begin
        cle.cl = inmsg.cl;
        cle.state = Dict_S;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_S;
        cle.perm = None;
        end

      end

      PutS: begin
        msg = fn_Resp(address,Put_Ack,cle.id,inmsg.src,cle.cl);
        send_fwd1 = tagged Valid msg;
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        if (fn_VectorCount (cle.sv) == 0) begin
        cle.state = Dict_I;
        cle.perm = None;

      end

        else begin
        cle.state = Dict_S;
        cle.perm = None;
        end

      end

      Upgrade: begin
        if (fn_IsElement (cle.sv,inmsg.src)) begin
        cle.sv = fn_RemoveElement(cle.sv,inmsg.src);
        msg = fn_RespAck(address,GetM_Ack_AD,cle.id,inmsg.src,cle.cl,fn_VectorCount (cle.sv));
        send_resp1 = tagged Valid msg;
        cle.state = Dict_M;
        cle.perm = None;
        msg = fn_Ack(address,Inv,inmsg.src,inmsg.src);
        send_multicast = tagged Valid tuple2(msg,cle.sv);
        cle.owner = inmsg.src;
        cle.sv = fn_Clear(cle.sv);

      end

        else begin
        msg = fn_RespAck(address,GetM_Ack_AD,cle.id,inmsg.src,cle.cl,fn_VectorCount (cle.sv));
        send_resp1 = tagged Valid msg;
        cle.state = Dict_M;
        cle.perm = None;
        msg = fn_Ack(address,Inv,inmsg.src,inmsg.src);
        send_multicast = tagged Valid tuple2(msg,cle.sv);
        cle.owner = inmsg.src;
        cle.sv = fn_Clear(cle.sv);
        end

      end

       default: stall = True;
    endcase
    end

endcase
return DictReturn { stall : stall, new_cle: cle, send_resp1: send_resp1, send_fwd1: send_fwd1, send_multicast: send_multicast};
endfunction


function Tuple2#(ENTRY_Cacheline_state#(w),Maybe#(Message#(a,w))) func_frm_core (ENTRY_Cacheline_state#(w) cle, Bit#(a) address, Access request);

  Message#(a,w) msg=unpack(0); 
  Maybe#(Message#(a,w)) send_req1 = tagged Invalid;

  if (cle.state == Cacheline_state_I && request == Load) begin
    msg = fn_Request(address,GetS,cle.id,tagged Directory);
    send_req1 = tagged Valid msg;
    cle.state = Cacheline_state_I_Load;
    cle.perm = None;
  end

  if (cle.state == Cacheline_state_I && request == Store) begin
    msg = fn_Request(address,GetM,cle.id,tagged Directory);
    send_req1 = tagged Valid msg;
    cle.acksReceived = 0;
    cle.state = Cacheline_state_I_Store;
    cle.perm = None;
  end


  if (cle.state == Cacheline_state_M && request == Evict) begin
    msg = fn_Resp(address,PutM,cle.id,tagged Directory,cle.cl);
    send_req1 = tagged Valid msg;
    cle.state = Cacheline_state_M_Evict;
    cle.perm = None;
  end

  if (cle.state == Cacheline_state_M && request == Load) begin
    cle.state = Cacheline_state_M;
    cle.perm = Store;
  end

  if (cle.state == Cacheline_state_M && request == Store) begin
    cle.state = Cacheline_state_M;
    cle.perm = Store;
  end


  if (cle.state == Cacheline_state_S && request == Evict) begin
    msg = fn_Request(address,PutS,cle.id,tagged Directory);
    send_req1 = tagged Valid msg;
    cle.state = Cacheline_state_S_Evict;
    cle.perm = None;
  end

  if (cle.state == Cacheline_state_S && request == Load) begin
    cle.state = Cacheline_state_S;
    cle.perm = Load;
  end

  if (cle.state == Cacheline_state_S && request == Store) begin
    msg = fn_Request(address,Upgrade,cle.id,tagged Directory);
    send_req1 = tagged Valid msg;
    cle.acksReceived = 0;
    cle.state = Cacheline_state_S_Store;
    cle.perm = Load;
  end


  return tuple2(cle, send_req1);

endfunction


endpackage