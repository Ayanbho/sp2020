package bridge_connectables;

	import axi4_axi4 ::*;
	import axi2axil ::*;
	import axi4lite_axi4lite ::*;
	import axi4lite_axi4 ::*;

	export axi4_axi4 ::*;
	export axi2axil ::*;
	export axi4lite_axi4lite ::*;
	export axi4lite_axi4 ::*;
	

endpackage
